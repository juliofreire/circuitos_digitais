library verilog;
use verilog.vl_types.all;
entity relatorio3_vlg_check_tst is
    port(
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end relatorio3_vlg_check_tst;
