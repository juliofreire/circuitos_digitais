library verilog;
use verilog.vl_types.all;
entity relatorio2_vlg_vec_tst is
end relatorio2_vlg_vec_tst;
