library verilog;
use verilog.vl_types.all;
entity relatorio3a is
    port(
        i0              : in     vl_logic;
        ia              : in     vl_logic;
        i2              : in     vl_logic;
        i3              : in     vl_logic;
        s0              : in     vl_logic;
        s1              : in     vl_logic;
        x               : out    vl_logic;
        x1              : out    vl_logic
    );
end relatorio3a;
