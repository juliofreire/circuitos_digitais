library verilog;
use verilog.vl_types.all;
entity relatorio3_vlg_sample_tst is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        i0              : in     vl_logic;
        i2              : in     vl_logic;
        i3              : in     vl_logic;
        ia              : in     vl_logic;
        s               : in     vl_logic;
        s0              : in     vl_logic;
        s1              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end relatorio3_vlg_sample_tst;
