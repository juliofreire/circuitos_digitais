library verilog;
use verilog.vl_types.all;
entity relatorio2_vlg_check_tst is
    port(
        s1              : in     vl_logic;
        s2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end relatorio2_vlg_check_tst;
