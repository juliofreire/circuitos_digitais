library verilog;
use verilog.vl_types.all;
entity relatorio5 is
    port(
        I3              : in     vl_logic;
        I2              : in     vl_logic;
        I1              : in     vl_logic;
        I0              : in     vl_logic;
        c               : in     vl_logic;
        Q3              : out    vl_logic;
        Q2              : out    vl_logic;
        Q1              : out    vl_logic;
        Q0              : out    vl_logic;
        O3              : out    vl_logic;
        O2              : out    vl_logic;
        O1              : out    vl_logic;
        O0              : out    vl_logic
    );
end relatorio5;
