library verilog;
use verilog.vl_types.all;
entity relatorio3a_vlg_vec_tst is
end relatorio3a_vlg_vec_tst;
