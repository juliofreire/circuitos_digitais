library verilog;
use verilog.vl_types.all;
entity projeto_final_vlg_check_tst is
    port(
        b1              : in     vl_logic;
        b2              : in     vl_logic;
        c0              : in     vl_logic;
        c1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end projeto_final_vlg_check_tst;
