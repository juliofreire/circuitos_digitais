library verilog;
use verilog.vl_types.all;
entity relatorio_vlg_vec_tst is
end relatorio_vlg_vec_tst;
