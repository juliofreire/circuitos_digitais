library verilog;
use verilog.vl_types.all;
entity relatorio3_vlg_vec_tst is
end relatorio3_vlg_vec_tst;
