library verilog;
use verilog.vl_types.all;
entity relatorio5_vlg_check_tst is
    port(
        O0              : in     vl_logic;
        O1              : in     vl_logic;
        O2              : in     vl_logic;
        O3              : in     vl_logic;
        Q0              : in     vl_logic;
        Q1              : in     vl_logic;
        Q2              : in     vl_logic;
        Q3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end relatorio5_vlg_check_tst;
