library verilog;
use verilog.vl_types.all;
entity relatorio5_vlg_vec_tst is
end relatorio5_vlg_vec_tst;
