library verilog;
use verilog.vl_types.all;
entity relatorio6_vlg_vec_tst is
end relatorio6_vlg_vec_tst;
