library verilog;
use verilog.vl_types.all;
entity relatorio_vlg_check_tst is
    port(
        a311            : in     vl_logic;
        a312            : in     vl_logic;
        a321            : in     vl_logic;
        a322            : in     vl_logic;
        c211            : in     vl_logic;
        c212            : in     vl_logic;
        c221            : in     vl_logic;
        c222            : in     vl_logic;
        d411            : in     vl_logic;
        d412            : in     vl_logic;
        d421            : in     vl_logic;
        d422            : in     vl_logic;
        id1             : in     vl_logic;
        id2             : in     vl_logic;
        id3             : in     vl_logic;
        q1              : in     vl_logic;
        q2              : in     vl_logic;
        ra31            : in     vl_logic;
        ra32            : in     vl_logic;
        rc21            : in     vl_logic;
        rc22            : in     vl_logic;
        rid1            : in     vl_logic;
        rid2            : in     vl_logic;
        rid3            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end relatorio_vlg_check_tst;
