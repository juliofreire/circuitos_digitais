library verilog;
use verilog.vl_types.all;
entity relatorio3a_vlg_check_tst is
    port(
        x               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end relatorio3a_vlg_check_tst;
