library verilog;
use verilog.vl_types.all;
entity relatorio3 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        s               : in     vl_logic;
        i0              : in     vl_logic;
        ia              : in     vl_logic;
        i2              : in     vl_logic;
        i3              : in     vl_logic;
        s0              : in     vl_logic;
        s1              : in     vl_logic;
        x1              : out    vl_logic;
        x2              : out    vl_logic;
        x3              : out    vl_logic
    );
end relatorio3;
